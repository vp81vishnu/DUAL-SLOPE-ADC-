* C:\Users\itops\Desktop\esim1\neww\neww.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/08/22 22:49:15

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_U5-Pad5_ Net-_U5-Pad6_ count24		
U7  Net-_U5-Pad6_ Net-_U5-Pad5_ Net-_U5-Pad4_ Net-_U5-Pad3_ Net-_U4-Pad~_ Net-_U3-Pad~_ Net-_U2-Pad~_ Net-_U1-Pad~_ adc_bridge_4		
v1  GND Net-_U5-Pad2_ DC		
v2  Net-_X1-Pad4_ GND DC		
v3  Net-_X1-Pad1_ GND DC		
v5  GND Net-_X1-Pad2_ DC		
U1  Net-_U1-Pad~_ plot_v1		
U2  Net-_U2-Pad~_ plot_v1		
U3  Net-_U3-Pad~_ plot_v1		
U4  Net-_U4-Pad~_ plot_v1		
U6  GND plot_v1		
U8  GND plot_v1		
X1  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_X1-Pad1_ Net-_X1-Pad4_ Net-_X1-Pad4_ GND avsd_opamp		
X2  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_X1-Pad1_ Net-_X1-Pad4_ Net-_U5-Pad1_ GND avsd_opamp		

.end
